library ieee;
use ieee.std_logic_1164.all;

entity REG_12 is
    port (
        clk : in std_logic;
        reset : in std_logic;
        enable : in std_logic;
        data_in : in std_logic_vector(11 downto 0);
        data_out : out std_logic_vector(11 downto 0)
    );
end entity REG_12;

architecture behavioral of REG_12 is
    signal reg : std_logic_vector(11 downto 0);
begin
    process(clk)
    begin
        if rising_edge(clk) then
            if reset = '1' then
                reg <= (others => '0');
            elsif enable = '1' then
                reg <= data_in;
            end if;
        end if;
    end process;

    data_out <= reg;
end architecture behavioral;